module selector(
    input wire a, b, select,
    output reg out
);
    
    assign out = in;
endmodule
