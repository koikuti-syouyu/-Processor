module template(
    input wire in,
    output reg out
);
    assign out = in;
endmodule
